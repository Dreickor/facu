library verilog;
use verilog.vl_types.all;
entity PARTED_vlg_vec_tst is
end PARTED_vlg_vec_tst;
