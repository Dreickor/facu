library verilog;
use verilog.vl_types.all;
entity sum_comp_vlg_vec_tst is
end sum_comp_vlg_vec_tst;
