-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 16 18:44:26 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PARTED IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        X : IN STD_LOGIC := '0';
        Led1 : OUT STD_LOGIC;
        Led2 : OUT STD_LOGIC;
        Led3 : OUT STD_LOGIC;
        Led4 : OUT STD_LOGIC
    );
END PARTED;

ARCHITECTURE BEHAVIOR OF PARTED IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state7,state6);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,X)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            Led1 <= '0';
            Led2 <= '0';
            Led3 <= '0';
            Led4 <= '0';
        ELSE
            Led1 <= '0';
            Led2 <= '0';
            Led3 <= '0';
            Led4 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((X = '1')) THEN
                        reg_fstate <= state6;
                    ELSIF ((X = '0')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    Led4 <= '0';

                    Led1 <= '0';

                    Led2 <= '0';

                    Led3 <= '0';
                WHEN state2 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    Led1 <= '0';
                    Led1 <= '1';
                    Led1 <= '1';
                    Led1 <= '0';
                WHEN state3 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state4;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    Led1 <= '1';
                    Led1 <= '1';
                    Led1 <= '1';
                    Led1 <= '1';
                WHEN state4 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    Led1 <= '0';
                    Led1 <= '0';
                    Led1 <= '1';

                    Led2 <= '1';
                WHEN state5 =>
                    IF ((X = '1')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    Led1 <= '1';
                    Led1 <= '0';
                    Led1 <= '0';
                    Led1 <= '0';
                WHEN state7 =>
                    IF ((X = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    Led1 <= '1';
                    Led1 <= '1';
                    Led1 <= '1';
                    Led1 <= '0';
                WHEN state6 =>
                    IF ((X = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    Led1 <= '0';
                    Led1 <= '0';

                    Led2 <= '1';

                    Led3 <= '1';
                WHEN OTHERS => 
                    Led1 <= 'X';
                    Led2 <= 'X';
                    Led3 <= 'X';
                    Led4 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
