library verilog;
use verilog.vl_types.all;
entity sum_comp_vlg_check_tst is
    port(
        ocout           : in     vl_logic;
        ores            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sum_comp_vlg_check_tst;
