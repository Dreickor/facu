library verilog;
use verilog.vl_types.all;
entity PARTEA_vlg_vec_tst is
end PARTEA_vlg_vec_tst;
