-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Nov 18 14:48:03 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Block2 IS 
	PORT
	(
		cin :  IN  STD_LOGIC;
		a0 :  IN  STD_LOGIC;
		a1 :  IN  STD_LOGIC;
		a2 :  IN  STD_LOGIC;
		a3 :  IN  STD_LOGIC;
		b0 :  IN  STD_LOGIC;
		b1 :  IN  STD_LOGIC;
		b2 :  IN  STD_LOGIC;
		b3 :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		res0 :  OUT  STD_LOGIC;
		res1 :  OUT  STD_LOGIC;
		res2 :  OUT  STD_LOGIC;
		res3 :  OUT  STD_LOGIC;
		cout :  OUT  STD_LOGIC;
		N :  OUT  STD_LOGIC;
		z :  OUT  STD_LOGIC;
		V :  OUT  STD_LOGIC
	);
END Block2;

ARCHITECTURE bdf_type OF Block2 IS 

COMPONENT partec
	PORT(a : IN STD_LOGIC;
		 b : IN STD_LOGIC;
		 cin : IN STD_LOGIC;
		 res : OUT STD_LOGIC;
		 cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	DFF_inst20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	DFF_inst21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	DFF_inst27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	DFF_inst19 :  STD_LOGIC;
SIGNAL	DFF_inst23 :  STD_LOGIC;
SIGNAL	DFF_inst28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	DFF_inst34 :  STD_LOGIC;


BEGIN 
res3 <= DFF_inst34;
N <= DFF_inst34;
SYNTHESIZED_WIRE_60 <= '1';
SYNTHESIZED_WIRE_61 <= '1';



b2v_inst : partec
PORT MAP(a => DFF_inst20,
		 b => SYNTHESIZED_WIRE_0,
		 cin => SYNTHESIZED_WIRE_56,
		 res => SYNTHESIZED_WIRE_62,
		 cout => SYNTHESIZED_WIRE_2);


b2v_inst1 : partec
PORT MAP(a => DFF_inst21,
		 b => SYNTHESIZED_WIRE_1,
		 cin => SYNTHESIZED_WIRE_2,
		 res => SYNTHESIZED_WIRE_64,
		 cout => SYNTHESIZED_WIRE_15);


SYNTHESIZED_WIRE_45 <= SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_5 AND SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_57;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_58);



SYNTHESIZED_WIRE_6 <= NOT(SYNTHESIZED_WIRE_59);



SYNTHESIZED_WIRE_8 <= NOT(SYNTHESIZED_WIRE_57);



PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_56 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_56 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_56 <= cin;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst19 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst19 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst19 <= b0;
END IF;
END PROCESS;


b2v_inst2 : partec
PORT MAP(a => DFF_inst27,
		 b => SYNTHESIZED_WIRE_14,
		 cin => SYNTHESIZED_WIRE_15,
		 res => SYNTHESIZED_WIRE_63,
		 cout => SYNTHESIZED_WIRE_40);


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst20 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst20 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst20 <= a0;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst21 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst21 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst21 <= a1;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_59 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_59 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_59 <= b3;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst23 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst23 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst23 <= b1;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_61,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	res0 <= '0';
ELSIF (SYNTHESIZED_WIRE_61 = '0') THEN
	res0 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	res0 <= SYNTHESIZED_WIRE_62;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_58 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	SYNTHESIZED_WIRE_58 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_58 <= a3;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_61,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	z <= '0';
ELSIF (SYNTHESIZED_WIRE_61 = '0') THEN
	z <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	z <= SYNTHESIZED_WIRE_30;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst27 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst27 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst27 <= a2;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_60,SYNTHESIZED_WIRE_60)
BEGIN
IF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst28 <= '0';
ELSIF (SYNTHESIZED_WIRE_60 = '0') THEN
	DFF_inst28 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst28 <= b2;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_61,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	res2 <= '0';
ELSIF (SYNTHESIZED_WIRE_61 = '0') THEN
	res2 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	res2 <= SYNTHESIZED_WIRE_63;
END IF;
END PROCESS;


b2v_inst3 : partec
PORT MAP(a => SYNTHESIZED_WIRE_58,
		 b => SYNTHESIZED_WIRE_39,
		 cin => SYNTHESIZED_WIRE_40,
		 res => SYNTHESIZED_WIRE_57,
		 cout => SYNTHESIZED_WIRE_51);


PROCESS(clk,SYNTHESIZED_WIRE_61,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	res1 <= '0';
ELSIF (SYNTHESIZED_WIRE_61 = '0') THEN
	res1 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	res1 <= SYNTHESIZED_WIRE_64;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_61,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	V <= '0';
ELSIF (SYNTHESIZED_WIRE_61 = '0') THEN
	V <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	V <= SYNTHESIZED_WIRE_45;
END IF;
END PROCESS;



PROCESS(clk,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	cout <= '0';
ELSIF (RISING_EDGE(clk)) THEN
	cout <= SYNTHESIZED_WIRE_48;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_61)
BEGIN
IF (SYNTHESIZED_WIRE_61 = '0') THEN
	DFF_inst34 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	DFF_inst34 <= SYNTHESIZED_WIRE_57;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_56 XOR DFF_inst19;


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_56 XOR DFF_inst23;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_56 XOR DFF_inst28;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_56 XOR SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_51 XOR SYNTHESIZED_WIRE_56;


SYNTHESIZED_WIRE_30 <= NOT(SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_62);


END bdf_type;